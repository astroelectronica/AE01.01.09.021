.title KiCad schematic
.include "models/C2012C0G2E102J085AA_p.mod"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/C2012X7R2E103K125AA_p.mod"
.include "models/C3216X5R1H106M160AB_p.mod"
.include "models/MAX4080T.FAM"
XU1 /VCC 0 C3216X5R1H106M160AB_p
XU2 /VCC 0 C2012X7R2A104K125AA_p
R1 /VIN /RSP 20
XU3 /RSP /RSN C2012C0G2E102J085AA_p
R4 /VOUT /RSN 20
R2 /VOUT /VIN 0.1
R3 /VOUT /VIN 0.1
XU4 /RSP /VCC NC_01 0 /VOCM NC_02 NC_03 /RSN MAX4080T
R5 /VOCM /CURRENT_FEEDBACK 100
XU5 /CURRENT_FEEDBACK 0 C2012X7R2E103K125AA_p
I1 /VOUT 0 {ILOAD}
V1 /VIN 0 {VSOURCE}
V2 /VCC 0 {VSUPPLY}
.end
